





//parameter WIDTH=8;
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//    FILE Name     :  d_flip_flop.sv                                                                             //
//                                                                                                                //
//    Description   :  D ff will trasfer the Data when Reset is low                                               //
//                                                                                                                //
//    Inputs        :  clk,reset,D                                                                                //
//                                                                                                                //
//    Outputs       :  Q                                                                                          //
//                                                                                                                //
                                                                                                                  //
//                                                                                                                //
//                                                                                                                //
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////










module d_flip_flop(
   input clk,
   input reset,
   input  D,
   output reg Q
   );

always@(posedge clk)
   
   begin
      if (reset) Q <=  0 ;
//      else if (D==1 || D ==0)  Q <=  D ;
      else Q<=D;
   end


endmodule

